----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:00:23 23.12.2012
-- Design Name: 
-- Module Name:    BatDecimator - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BatDecimator is
	Port (
		i_DC_RESET						: in  STD_LOGIC;
		i_DC_USRCLK						: in  STD_LOGIC;								-- User clock 100 MHz
		
		i_DC_625KHZ						: in  STD_LOGIC;								-- 0: 312500 1: 625 KHZ
				
		i_DC_DataAv						: in  STD_LOGIC;								-- new data available in DataIn
		i_DC_DataAvOut					: out STD_LOGIC;								-- new data available generated by decimator
		
		i_DC_R_DataIn					: in  std_logic_vector(23 downto 0);	-- new data from ADC
		i_DC_L_DataIn					: in  std_logic_vector(23 downto 0);	-- new data from ADC
		i_DC_R_DataOut					: out std_logic_vector(23 downto 0);	-- data for DAC
		i_DC_L_DataOut					: out std_logic_vector(23 downto 0);	-- data for DAC
		i_DC_Random                : in	std_logic_vector(31 downto 0)		-- Random data	
	);
end BatDecimator;

--##################################################################################
--#	Architecture
--#
--#
--##################################################################################
architecture Behavioral of BatDecimator is
--##################################################################################
--#	Constants
--#
--#
--##################################################################################


--##################################################################################
--#	Components
--#
--#
--##################################################################################

component Decimator
	port (
		clk								: in std_logic;
		ce									: in std_logic;
		nd									: in std_logic;
		rfd								: out std_logic;
		rdy								: out std_logic;
		chan_in							: out std_logic_vector(0 downto 0);
		chan_out							: out std_logic_vector(0 downto 0);
		din								: in std_logic_vector(23 downto 0);
		dout								: out std_logic_vector(49 downto 0));
end component;

component BatDither
	generic(
		dBits								: integer;
		qBits								: integer;
		ditherBits						: integer										-- min ((dBits-qBits) + 1)
	);

   port (
		clk								: in std_logic;
		nd									: in std_logic;
		bypass							: in std_logic;

		dither							: in signed(ditherBits-1 downto 0);
		d									: in signed(dBits-1 downto 0);
		q									: out std_logic_vector(qBits-1 downto 0)
	);
end component;

--##################################################################################
--#	Signals
--#
--#
--##################################################################################
-----------------------
-- Decimator divider --
-----------------------
signal	s_FilterIn						: signed(23 downto 0);					-- the filter input
signal	s_DC_Out							: std_logic_vector(49 downto 0) := (others => '0');	-- of filtering
signal	s_DC_OutDith					: std_logic_vector(23 downto 0) := (others => '0');	-- dithered version of filtering
signal	s_DC_OutReg						: std_logic_vector(23 downto 0) := (others => '0');	-- save result of first channel until second channel is ready

signal	s_FilterRdy						: std_logic := '0';						-- new outputdata availabe at filter
signal	s_RdyForData					: std_logic := '0';						-- Filter is ready to accept new data
signal	s_EN								: std_logic := '0';						-- Enable signal for Multiplier and Filter (to save a bit of power)
signal	s_ChanIn							: std_logic_vector(0 downto 0) := "0";		-- Input channel selector
signal	s_ChanOut						: std_logic_vector(0 downto 0) := "0";		-- Output channel selector
signal	s_ND								: std_logic := '0';						-- New Data signal
signal	s_DithNd							: std_logic := '0';						-- new dither data

signal	s_DithIn							: signed(47 downto 0);					-- the dither input


-- DC Read Statemachine states
TYPE 		RSTATE_TYPE IS (St_R0, St_R1, St_R2, St_R3, St_R4, St_R5);
signal 	s_RState							: RSTATE_TYPE := St_R0;
-- DC Feed Statemachine states
TYPE 		FSTATE_TYPE IS (St_F0, St_F1, St_F2, St_F3);
signal 	s_FState							: FSTATE_TYPE := St_F0;

--##################################################################################
--#	Architecture Body
--#
--#
--##################################################################################
begin

inst_Decimator: Decimator
	port map (
		clk 								=> i_DC_USRCLK,
		ce 								=> s_EN,
		nd 								=> s_ND,
		chan_in 							=> s_ChanIn,
		chan_out 						=> s_ChanOut,
		rfd 								=> s_RdyForData,
		rdy 								=> s_FilterRdy,
		din 								=> std_logic_vector(s_FilterIn),
		dout 								=> s_DC_Out
	);
	
inst_DecDither: BatDither
	generic map(
		dBits								=> 48,
		qBits								=> 24,
		ditherBits						=> 25										-- min ((dBits-qBits) + 1)
	)
 	port map (
		clk								=> i_DC_USRCLK,
		nd									=> s_DithNd,
		bypass							=> '0',

		dither							=> signed(i_DC_Random(24 downto 0)),
		d									=> s_DithIn,
		q									=> s_DC_OutDith
	);

s_DithIn <= signed(s_DC_Out(49) & s_DC_Out(46 downto 0));

-----------------------------------------------------------
-- Feed Decimator Filter
-----------------------------------------------------------
DecFeedFIRProc: process(i_DC_USRCLK)
begin
	if rising_edge(i_DC_USRCLK) then
		-- Reset
		if i_DC_RESET = '1' then
			s_EN <= '0';
			s_ND <= '0';
			s_FilterIn <= (others => '0');
		else
		-- Clock
			s_ND <= '0';																	-- reset ND signal
			s_EN <= '1';
			case s_FState is
				when St_F0 =>
					if i_DC_DataAv = '1' and s_ChanIn = "0" then					-- new data available, sync on channel 0
						s_FState <= St_F1;                                 	-- next state
					else
						s_FState <= St_F0;                                 	-- keep state
					end if;
				when St_F1 =>
					if s_RdyForData = '1' then											-- Filter ready to accept data?
						s_FilterIn <= signed(i_DC_R_DataIn);						-- feed with right channel
						s_ND <= '1';														-- take over data to filter
						s_FState <= St_F2;                                 	-- next state
					else
						s_FState <= St_F1;                                 	-- keep state
					end if;
				when St_F2 =>
						s_FState <= St_F3;                                 	-- next state
				when St_F3 =>
					if s_RdyForData = '1' and s_ChanIn = "1" then				-- Filter ready to accept data?
						s_FilterIn <= signed(i_DC_L_DataIn);						-- feed with left channel
						s_ND <= '1';														-- take over data to filter
						s_FState <= St_F0;                                 	-- default state
					else
						s_FState <= St_F3;                                 	-- keep state
					end if;
			end case;
		end if;
	end if;
end process DecFeedFIRProc;

-----------------------------------------------------------
-- Write result
-----------------------------------------------------------
DecOutProc: process(i_DC_USRCLK)
begin
	if rising_edge(i_DC_USRCLK) then
		-- Reset
		if i_DC_RESET = '1' then
			i_DC_R_DataOut <= (others => '0');										-- reset value for output signal
			i_DC_L_DataOut <= (others => '0');										-- reset value for output signal
			s_RState <= St_R0;
			s_DithNd <= '0';
			i_DC_DataAvOut <= '0';
		else
		-- Clock
		   if i_DC_625KHZ = '1' then
				s_DithNd <= '0';															-- reset DithND every clock			
				i_DC_DataAvOut <= '0';
				case s_RState is
					when St_R0 =>
						if s_FilterRdy = '1' and s_ChanOut = "0" then			-- now we have the filtered value in s_FilterOut, sync on channel 0
							s_DithNd <= '1';
							s_RState <= St_R1;											-- next state
						else
							s_RState <= St_R0;                                	-- keep state
						end if;
					when St_R1 =>															-- wait one cycle to be sure to have dithered data
						s_RState <= St_R2;												-- next state
					when St_R2 =>															-- here we should have dithered data available
						s_DC_OutReg <= s_DC_OutDith;									-- right channel ready
						s_RState <= St_R3;												-- next state
					when St_R3 =>															-- wait for Filter ready to disappear
						if s_FilterRdy = '1' then										-- this can only be channel 1
							s_DithNd <= '1';
							s_RState <= St_R4;											-- next state
						else
							s_RState <= St_R3;                                	-- keep state
						end if;
					when St_R4 =>															-- wait one cycle to be sure to have dithered data
						s_RState <= St_R5;												-- next state
					when St_R5 =>															-- wait for Filter ready to diappear
						i_DC_L_DataOut <= s_DC_OutDith;								-- left channel ready
						i_DC_R_DataOut <= s_DC_OutReg;								-- change both channels at the same time
						i_DC_DataAvOut <= '1';
						s_RState <= St_R0;												-- next state
				end case;
			else																				-- we are in 3125.5 KHZ mode, do nothing
				i_DC_DataAvOut <= i_DC_DataAv;
				i_DC_R_DataOut <= i_DC_R_DataIn;
				i_DC_L_DataOut <= i_DC_L_DataIn;
			end if;
		end if;
	end if;
end process DecOutProc;

end Behavioral;